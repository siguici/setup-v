module main

fn test_welcome() {
	assert welcome('Sigui') == 'Hello, Sigui. Welcome to V!'
}
